.SUBCKT PORT_1 NODE_TOP NODE_BOT
R0 NODE_TOP NODE_MID [1552.44605269    0.            0.            0.            0.
    0.            0.            0.            0.            0.
    0.            0.            0.            0.            0.        ]
L0 NODE_MID NODE_BOT [0.00023583 0.         0.         0.         0.         0.
 0.         0.         0.         0.         0.         0.
 0.         0.         0.        ]
RA1 NODE_TOP NODE_12 2489.4544755897487
RB1 NODE_13 NODE_BOT 29193.0421254109
L1 NODE_12 NODE_13 0.01400149301402511
C1 NODE_13 NODE_BOT 1.8900814584037922e-10
RA2 NODE_TOP NODE_22 2489.4544755897487
RB2 NODE_23 NODE_BOT 29193.0421254109
L2 NODE_22 NODE_23 0.01400149301402511
C2 NODE_23 NODE_BOT 1.8900814584037922e-10
RA3 NODE_TOP NODE_32 2342.6087550552575
RB3 NODE_33 NODE_BOT 19725.31065182912
L3 NODE_32 NODE_33 0.014946130148356935
C3 NODE_33 NODE_BOT 3.1752520448264074e-10
RA4 NODE_TOP NODE_42 2342.6087550552575
RB4 NODE_43 NODE_BOT 19725.31065182912
L4 NODE_42 NODE_43 0.014946130148356935
C4 NODE_43 NODE_BOT 3.1752520448264074e-10
RA5 NODE_TOP NODE_52 1227.3046700546643
RB5 NODE_53 NODE_BOT 3649.7989824657466
L5 NODE_52 NODE_53 0.046990577062158666
C5 NODE_53 NODE_BOT 1.149011232182718e-08
RA6 NODE_TOP NODE_62 1227.3046700546643
RB6 NODE_63 NODE_BOT 3649.7989824657466
L6 NODE_62 NODE_63 0.046990577062158666
C6 NODE_63 NODE_BOT 1.149011232182718e-08
RA7 NODE_TOP NODE_72 2328.269746868149
RB7 NODE_73 NODE_BOT 9055.704167097294
L7 NODE_72 NODE_73 0.014522386787622006
C7 NODE_73 NODE_BOT 6.802795124193373e-10
RA8 NODE_TOP NODE_82 2328.269746868149
RB8 NODE_83 NODE_BOT 9055.704167097294
L8 NODE_82 NODE_83 0.014522386787622006
C8 NODE_83 NODE_BOT 6.802795124193373e-10
RA9 NODE_TOP NODE_92 504.81132026190807
RB9 NODE_93 NODE_BOT 8351.56233120223
L9 NODE_92 NODE_93 0.010333235623323169
C9 NODE_93 NODE_BOT 2.38198505133009e-09
RA10 NODE_TOP NODE_102 504.81132026190807
RB10 NODE_103 NODE_BOT 8351.56233120223
L10 NODE_102 NODE_103 0.010333235623323169
C10 NODE_103 NODE_BOT 2.38198505133009e-09
RA11 NODE_TOP NODE_112 105.7490398791496
RB11 NODE_113 NODE_BOT 12801.351557040567
L11 NODE_112 NODE_113 0.010302480869210389
C11 NODE_113 NODE_BOT 7.001699585102146e-09
RA12 NODE_TOP NODE_122 105.7490398791496
RB12 NODE_123 NODE_BOT 12801.351557040567
L12 NODE_122 NODE_123 0.010302480869210389
C12 NODE_123 NODE_BOT 7.001699585102146e-09
RA13 NODE_TOP NODE_132 13.093212299901783
RB13 NODE_133 NODE_BOT 32695.042324284084
L13 NODE_132 NODE_133 0.01416476077462686
C13 NODE_133 NODE_BOT 4.623178540795888e-08
RA14 NODE_TOP NODE_142 13.093212299901783
RB14 NODE_143 NODE_BOT 32695.042324284084
L14 NODE_142 NODE_143 0.01416476077462686
C14 NODE_143 NODE_BOT 4.623178540795888e-08
.ENDS PORT_1

.SUBCKT PORT_2 NODE_TOP NODE_BOT
R0 NODE_TOP NODE_MID [1552.44605269    0.            0.            0.            0.
    0.            0.            0.            0.            0.
    0.            0.            0.            0.            0.        ]
L0 NODE_MID NODE_BOT [0.00023583 0.         0.         0.         0.         0.
 0.         0.         0.         0.         0.         0.
 0.         0.         0.        ]
RA1 NODE_TOP NODE_12 1323.191138540788
RB1 NODE_13 NODE_BOT 18295.054780375176
L1 NODE_12 NODE_13 0.007976542976268496
C1 NODE_13 NODE_BOT 3.36469513939152e-10
RA2 NODE_TOP NODE_22 1323.191138540788
RB2 NODE_23 NODE_BOT 18295.054780375176
L2 NODE_22 NODE_23 0.007976542976268496
C2 NODE_23 NODE_BOT 3.36469513939152e-10
RA3 NODE_TOP NODE_32 1234.5126407232858
RB3 NODE_33 NODE_BOT 13675.002293257381
L3 NODE_32 NODE_33 0.008996967202410664
C3 NODE_33 NODE_BOT 5.445370854671201e-10
RA4 NODE_TOP NODE_42 1234.5126407232858
RB4 NODE_43 NODE_BOT 13675.002293257381
L4 NODE_42 NODE_43 0.008996967202410664
C4 NODE_43 NODE_BOT 5.445370854671201e-10
RA5 NODE_TOP NODE_52 721.5317214244827
RB5 NODE_53 NODE_BOT 5286.330743698678
L5 NODE_52 NODE_53 0.04771404729865732
C5 NODE_53 NODE_BOT 1.4721847176444464e-08
RA6 NODE_TOP NODE_62 721.5317214244827
RB6 NODE_63 NODE_BOT 5286.330743698678
L6 NODE_62 NODE_63 0.04771404729865732
C6 NODE_63 NODE_BOT 1.4721847176444464e-08
RA7 NODE_TOP NODE_72 280.40150214518553
RB7 NODE_73 NODE_BOT 15184.32804213757
L7 NODE_72 NODE_73 0.00725890692076973
C7 NODE_73 NODE_BOT 1.798175354108358e-09
RA8 NODE_TOP NODE_82 280.40150214518553
RB8 NODE_83 NODE_BOT 15184.32804213757
L8 NODE_82 NODE_83 0.00725890692076973
C8 NODE_83 NODE_BOT 1.798175354108358e-09
RA9 NODE_TOP NODE_92 876.8876637449885
RB9 NODE_93 NODE_BOT 8640.137743050336
L9 NODE_92 NODE_93 0.013211162611109512
C9 NODE_93 NODE_BOT 1.7817020963983593e-09
RA10 NODE_TOP NODE_102 876.8876637449885
RB10 NODE_103 NODE_BOT 8640.137743050336
L10 NODE_102 NODE_103 0.013211162611109512
C10 NODE_103 NODE_BOT 1.7817020963983593e-09
RA11 NODE_TOP NODE_112 51.14102974085793
RB11 NODE_113 NODE_BOT 39701.37535748197
L11 NODE_112 NODE_113 0.010925699831762859
C11 NODE_113 NODE_BOT 6.6487306441183685e-09
RA12 NODE_TOP NODE_122 51.14102974085793
RB12 NODE_123 NODE_BOT 39701.37535748197
L12 NODE_122 NODE_123 0.010925699831762859
C12 NODE_123 NODE_BOT 6.6487306441183685e-09
RA13 NODE_TOP NODE_132 37.80461911681765
RB13 NODE_133 NODE_BOT 5303.533341089189
L13 NODE_132 NODE_133 0.010975670801268617
C13 NODE_133 NODE_BOT 5.9263318954424074e-08
RA14 NODE_TOP NODE_142 37.80461911681765
RB14 NODE_143 NODE_BOT 5303.533341089189
L14 NODE_142 NODE_143 0.010975670801268617
C14 NODE_143 NODE_BOT 5.9263318954424074e-08
.ENDS PORT_2

.SUBCKT PORT_3 NODE_TOP NODE_BOT
R0 NODE_TOP NODE_MID [1552.44605269    0.            0.            0.            0.
    0.            0.            0.            0.            0.
    0.            0.            0.            0.            0.        ]
L0 NODE_MID NODE_BOT [0.00023583 0.         0.         0.         0.         0.
 0.         0.         0.         0.         0.         0.
 0.         0.         0.        ]
RA1 NODE_TOP NODE_12 2489.4544755894785
RB1 NODE_13 NODE_BOT 29193.042125412358
L1 NODE_12 NODE_13 0.014001493014024815
C1 NODE_13 NODE_BOT 1.8900814584038602e-10
RA2 NODE_TOP NODE_22 2489.4544755894785
RB2 NODE_23 NODE_BOT 29193.042125412358
L2 NODE_22 NODE_23 0.014001493014024815
C2 NODE_23 NODE_BOT 1.8900814584038602e-10
RA3 NODE_TOP NODE_32 2342.6087550546313
RB3 NODE_33 NODE_BOT 19725.310651831835
L3 NODE_32 NODE_33 0.014946130148356402
C3 NODE_33 NODE_BOT 3.1752520448266944e-10
RA4 NODE_TOP NODE_42 2342.6087550546313
RB4 NODE_43 NODE_BOT 19725.310651831835
L4 NODE_42 NODE_43 0.014946130148356402
C4 NODE_43 NODE_BOT 3.1752520448266944e-10
RA5 NODE_TOP NODE_52 1227.3046700546108
RB5 NODE_53 NODE_BOT 3649.7989824657243
L5 NODE_52 NODE_53 0.04699057706215789
C5 NODE_53 NODE_BOT 1.1490112321827589e-08
RA6 NODE_TOP NODE_62 1227.3046700546108
RB6 NODE_63 NODE_BOT 3649.7989824657243
L6 NODE_62 NODE_63 0.04699057706215789
C6 NODE_63 NODE_BOT 1.1490112321827589e-08
RA7 NODE_TOP NODE_72 2328.269746867675
RB7 NODE_73 NODE_BOT 9055.704167097623
L7 NODE_72 NODE_73 0.014522386787621409
C7 NODE_73 NODE_BOT 6.802795124194218e-10
RA8 NODE_TOP NODE_82 2328.269746867675
RB8 NODE_83 NODE_BOT 9055.704167097623
L8 NODE_82 NODE_83 0.014522386787621409
C8 NODE_83 NODE_BOT 6.802795124194218e-10
RA9 NODE_TOP NODE_92 504.8113202619061
RB9 NODE_93 NODE_BOT 8351.562331202555
L9 NODE_92 NODE_93 0.010333235623323365
C9 NODE_93 NODE_BOT 2.3819850513300506e-09
RA10 NODE_TOP NODE_102 504.8113202619061
RB10 NODE_103 NODE_BOT 8351.562331202555
L10 NODE_102 NODE_103 0.010333235623323365
C10 NODE_103 NODE_BOT 2.3819850513300506e-09
RA11 NODE_TOP NODE_112 105.74903987914725
RB11 NODE_113 NODE_BOT 12801.351557041327
L11 NODE_112 NODE_113 0.010302480869210602
C11 NODE_113 NODE_BOT 7.001699585102007e-09
RA12 NODE_TOP NODE_122 105.74903987914725
RB12 NODE_123 NODE_BOT 12801.351557041327
L12 NODE_122 NODE_123 0.010302480869210602
C12 NODE_123 NODE_BOT 7.001699585102007e-09
RA13 NODE_TOP NODE_132 13.09321229990291
RB13 NODE_133 NODE_BOT 32695.04232428017
L13 NODE_132 NODE_133 0.014164760774626863
C13 NODE_133 NODE_BOT 4.623178540795887e-08
RA14 NODE_TOP NODE_142 13.09321229990291
RB14 NODE_143 NODE_BOT 32695.04232428017
L14 NODE_142 NODE_143 0.014164760774626863
C14 NODE_143 NODE_BOT 4.623178540795887e-08
.ENDS PORT_3

.END