.SUBCKT PORT_0 NODE_TOP NODE_BOT
RA0 NODE_TOP NODE_02 14004.992867332383
RB0 NODE_03 NODE_BOT 0.0
L0 NODE_02 NODE_03 2228.9586305278176
C0 NODE_03 NODE_BOT 0.0
RA1 NODE_TOP NODE_12 -2446.054538269003
RB1 NODE_13 NODE_BOT 0.0
L1 NODE_12 NODE_13 -131.73494928204454
C1 NODE_13 NODE_BOT 0.0
RA2 NODE_TOP NODE_22 977.1927139139752
RB2 NODE_23 NODE_BOT 0.0
L2 NODE_22 NODE_23 30.61380682687892
C2 NODE_23 NODE_BOT 0.0
RA3 NODE_TOP NODE_32 -690.0528169014085
RB3 NODE_33 NODE_BOT 0.0
L3 NODE_32 NODE_33 -12.575452716297788
C3 NODE_33 NODE_BOT 0.0
RA4 NODE_TOP NODE_42 774.0214983178796
RB4 NODE_43 NODE_BOT 0.0
L4 NODE_42 NODE_43 8.205464839583161
C4 NODE_43 NODE_BOT 0.0
RA5 NODE_TOP NODE_52 -1694.1963119678212
RB5 NODE_53 NODE_BOT 0.0
L5 NODE_52 NODE_53 -10.44768322624458
C5 NODE_53 NODE_BOT 0.0
RA6 NODE_TOP NODE_62 1093.2375449008277
RB6 NODE_63 NODE_BOT 0.0
L6 NODE_62 NODE_63 0.5205893070956322
C6 NODE_63 NODE_BOT 0.0
RA7 NODE_TOP NODE_72 1.032015411430144
RB7 NODE_73 NODE_BOT 0.0
L7 NODE_72 NODE_73 0.00022933675809558757
C7 NODE_73 NODE_BOT 0.0
RA8 NODE_TOP NODE_82 -1.3434236186348862
RB8 NODE_83 NODE_BOT 0.0
L8 NODE_82 NODE_83 -0.00021668472372697725
C8 NODE_83 NODE_BOT 0.0
RA9 NODE_TOP NODE_92 1.350938136592688
RB9 NODE_93 NODE_BOT 0.0
L9 NODE_92 NODE_93 0.00021443122118580465
C9 NODE_93 NODE_BOT 0.0
RA10 NODE_TOP NODE_102 -0.23681502890173411
RB10 NODE_103 NODE_BOT 0.0
L10 NODE_102 NODE_103 -5.780346820809249e-06
C10 NODE_103 NODE_BOT 0.0
RA11 NODE_TOP NODE_112 0.1414951768488746
RB11 NODE_113 NODE_BOT 0.0
L11 NODE_112 NODE_113 3.215434083601286e-06
C11 NODE_113 NODE_BOT 0.0
RA12 NODE_TOP NODE_122 -0.29835911602209947
RB12 NODE_123 NODE_BOT 0.0
L12 NODE_122 NODE_123 -5.524861878453038e-06
C12 NODE_123 NODE_BOT 0.0
RA13 NODE_TOP NODE_132 1.1837324199327577
RB13 NODE_133 NODE_BOT 0.0
L13 NODE_132 NODE_133 1.5784572159171624e-05
C13 NODE_133 NODE_BOT 0.0
RA14 NODE_TOP NODE_142 -1807115.6428894137
RB14 NODE_143 NODE_BOT 1807116.142903765
L14 NODE_142 NODE_143 0.13579576317218903
C14 NODE_143 NODE_BOT 4.1582814907654096e-14
RA15 NODE_TOP NODE_152 -1807115.6428894137
RB15 NODE_153 NODE_BOT 1807116.142903765
L15 NODE_152 NODE_153 0.13579576317218903
C15 NODE_153 NODE_BOT 4.1582814907654096e-14
RA16 NODE_TOP NODE_162 -9518.73669634292
RB16 NODE_163 NODE_BOT 9519.336691757899
L16 NODE_162 NODE_163 0.004198505332101771
C16 NODE_163 NODE_BOT 4.633412640059169e-11
RA17 NODE_TOP NODE_172 -9518.73669634292
RB17 NODE_173 NODE_BOT 9519.336691757899
L17 NODE_172 NODE_173 0.004198505332101771
C17 NODE_173 NODE_BOT 4.633412640059169e-11
.PLOT AC VM(NODE_TOP)
.ENDS PORT_0

.END